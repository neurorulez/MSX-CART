--
--  vga.vhd
--   VGA up-scan converter.
--
--  Copyright (C) 2006 Kunihiko Ohnaka
--  All rights reserved.
--                                     http://www.ohnaka.jp/ese-vdp/
--
--  –{ƒ\ƒtƒgƒEƒFƒA‚¨‚æ‚Ñ–{ƒ\ƒtƒgƒEƒFƒA‚ÉŠî‚Ã‚¢‚Äì¬‚³‚ê‚½”h¶•¨‚ÍAˆÈ‰º‚ÌðŒ‚ð
--  –ž‚½‚·ê‡‚ÉŒÀ‚èAÄ”Ð•z‚¨‚æ‚ÑŽg—p‚ª‹–‰Â‚³‚ê‚Ü‚·B
--
--  1.ƒ\[ƒXƒR[ƒhŒ`Ž®‚ÅÄ”Ð•z‚·‚éê‡Aã‹L‚Ì’˜ìŒ •\Ž¦A–{ðŒˆê——A‚¨‚æ‚Ñ‰º‹L
--    –ÆÓð€‚ð‚»‚Ì‚Ü‚Ü‚ÌŒ`‚Å•ÛŽ‚·‚é‚±‚ÆB
--  2.ƒoƒCƒiƒŠŒ`Ž®‚ÅÄ”Ð•z‚·‚éê‡A”Ð•z•¨‚É•t‘®‚ÌƒhƒLƒ…ƒƒ“ƒg“™‚ÌŽ‘—¿‚ÉAã‹L‚Ì
--    ’˜ìŒ •\Ž¦A–{ðŒˆê——A‚¨‚æ‚Ñ‰º‹L–ÆÓð€‚ðŠÜ‚ß‚é‚±‚ÆB
--  3.‘–Ê‚É‚æ‚éŽ–‘O‚Ì‹–‰Â‚È‚µ‚ÉA–{ƒ\ƒtƒgƒEƒFƒA‚ð”Ì”„A‚¨‚æ‚Ñ¤‹Æ“I‚È»•i‚âŠˆ“®
--    ‚ÉŽg—p‚µ‚È‚¢‚±‚ÆB
--
--  –{ƒ\ƒtƒgƒEƒFƒA‚ÍA’˜ìŒ ŽÒ‚É‚æ‚Á‚ÄuŒ»ó‚Ì‚Ü‚Üv’ñ‹Ÿ‚³‚ê‚Ä‚¢‚Ü‚·B’˜ìŒ ŽÒ‚ÍA
--  “Á’è–Ú“I‚Ö‚Ì“K‡«‚Ì•ÛØA¤•i«‚Ì•ÛØA‚Ü‚½‚»‚ê‚ÉŒÀ’è‚³‚ê‚È‚¢A‚¢‚©‚È‚é–¾Ž¦
--  “I‚à‚µ‚­‚ÍˆÃ–Ù‚È•ÛØÓ”C‚à•‰‚¢‚Ü‚¹‚ñB’˜ìŒ ŽÒ‚ÍAŽ–—R‚Ì‚¢‚©‚ñ‚ð–â‚í‚¸A‘¹ŠQ
--  ”­¶‚ÌŒ´ˆö‚¢‚©‚ñ‚ð–â‚í‚¸A‚©‚ÂÓ”C‚Ìª‹’‚ªŒ_–ñ‚Å‚ ‚é‚©ŒµŠiÓ”C‚Å‚ ‚é‚©i‰ßŽ¸
--  ‚»‚Ì‘¼‚Ìj•s–@sˆ×‚Å‚ ‚é‚©‚ð–â‚í‚¸A‰¼‚É‚»‚Ì‚æ‚¤‚È‘¹ŠQ‚ª”­¶‚·‚é‰Â”\«‚ð’m‚ç
--  ‚³‚ê‚Ä‚¢‚½‚Æ‚µ‚Ä‚àA–{ƒ\ƒtƒgƒEƒFƒA‚ÌŽg—p‚É‚æ‚Á‚Ä”­¶‚µ‚½i‘ã‘Ö•i‚Ü‚½‚Í‘ã—pƒT
--  [ƒrƒX‚Ì’²’BAŽg—p‚Ì‘rŽ¸Aƒf[ƒ^‚Ì‘rŽ¸A—˜‰v‚Ì‘rŽ¸A‹Æ–±‚Ì’†’f‚àŠÜ‚ßA‚Ü‚½‚»
--  ‚ê‚ÉŒÀ’è‚³‚ê‚È‚¢j’¼Ú‘¹ŠQAŠÔÚ‘¹ŠQA‹ô”­“I‚È‘¹ŠQA“Á•Ê‘¹ŠQA’¦”±“I‘¹ŠQA‚Ü
--  ‚½‚ÍŒ‹‰Ê‘¹ŠQ‚É‚Â‚¢‚ÄAˆêØÓ”C‚ð•‰‚í‚È‚¢‚à‚Ì‚Æ‚µ‚Ü‚·B
--
--  Note that above Japanese version license is the formal document.
--  The following translation is only for reference.
--
--  Redistribution and use of this software or any derivative works,
--  are permitted provided that the following conditions are met:
--
--  1. Redistributions of source code must retain the above copyright
--     notice, this list of conditions and the following disclaimer.
--  2. Redistributions in binary form must reproduce the above
--     copyright notice, this list of conditions and the following
--     disclaimer in the documentation and/or other materials
--     provided with the distribution.
--  3. Redistributions may not be sold, nor may they be used in a 
--     commercial product or activity without specific prior written
--     permission.
--
--  THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS 
--  "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT 
--  LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS
--  FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
--  COPYRIGHT OWNER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT,
--  INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING,
--  BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
--  LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER 
--  CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT
--  LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN
--  ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
--  POSSIBILITY OF SUCH DAMAGE.
--
-------------------------------------------------------------------------------
-- Memo
--   Japanese comment lines are starts with "JP:".
--   JP: “ú–{Œê‚ÌƒRƒƒ“ƒgs‚Í JP:‚ð“ª‚É•t‚¯‚éŽ–‚É‚·‚é
--
-------------------------------------------------------------------------------
-- Revision History
--
-- 29th,October,2006 modified by Kunihiko Ohnaka
--   - Insert the license text.
--   - Add the document part below.
--
-- ?th,August,2006 modified by Kunihiko Ohnaka
--   - Move the equalization pulse generator from
--     vdp.vhd.
--
-- 20th,August,2006 modified by Kunihiko Ohnaka
--  - Change field mapping algorithm when interlace
--    mode is enabled.
--        even field  -> even line (odd  line is blacK)
--        odd  field  -> odd line  (even line is blacK)
--
-- 13th,October,2003 created by Kunihiko Ohnaka
-- JP: VDP‚ÌƒRƒA‚ÌŽÀ‘•‚Æ•\Ž¦ƒfƒoƒCƒX‚Ö‚Ìo—Í‚ð•Êƒ\[ƒX‚É‚µ‚½D
-- TRANSLATED: Implemented VDP core and output to display device as separate sources.
--
-------------------------------------------------------------------------------
-- Document
--
-- JP: ESE-VDPƒRƒA(vdp.vhd)‚ª¶¬‚µ‚½ƒrƒfƒIM†‚ðAVGAƒ^ƒCƒ~ƒ“ƒO‚É
-- JP: •ÏŠ·‚·‚éƒAƒbƒvƒXƒLƒƒƒ“ƒRƒ“ƒo[ƒ^‚Å‚·B
-- JP: NTSC‚Í…•½“¯ŠúŽü”g”‚ª15.7KHzA‚’¼“¯ŠúŽü”g”‚ª60Hz‚Å‚·‚ªA
-- JP: VGA‚Ì…•½“¯ŠúŽü”g”‚Í31.5KHzA‚’¼“¯ŠúŽü”g”‚Í60Hz‚Å‚ ‚èA
-- JP: ƒ‰ƒCƒ“”‚¾‚¯‚ª‚Ù‚Ú”{‚É‚È‚Á‚½‚æ‚¤‚Èƒ^ƒCƒ~ƒ“ƒO‚É‚È‚è‚Ü‚·B
-- JP: ‚»‚±‚ÅAvdp‚ð ntscƒ‚[ƒh‚Å“®‚©‚µAŠeƒ‰ƒCƒ“‚ð”{‚Ì‘¬“x‚Å
-- JP: “ñ“x•`‰æ‚·‚é‚±‚Æ‚ÅƒXƒLƒƒƒ“ƒRƒ“ƒo[ƒg‚ðŽÀŒ»‚µ‚Ä‚¢‚Ü‚·B
--
-- TRANSLATION BY GOOGLE
-- JP: Video signal generated by ESE-VDP core (vdp.vhd) to VGA timing
-- JP: Up scan converter to convert.
-- JP: NTSC has a horizontal sync frequency of 15.7 KHz and a vertical sync frequency of 60 Hz.
-- JP: VGA horizontal sync frequency is 31.5 KHz, vertical sync frequency is 60 Hz,
-- JP: Timing is almost doubled only by the number of lines.
-- JP: So, move vdp in ntsc mode and double each speed
-- JP: Scan conversion is realized by drawing twice.
--

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use work.vdp_package.all;

entity vdp_vga is
  port(
    -- VDP clock ... 21.477MHz
    clk21m  : in std_logic;
    reset   : in std_logic;

    -- Video Input
    videoRin : in std_logic_vector( 5 downto 0);
    videoGin : in std_logic_vector( 5 downto 0);
    videoBin : in std_logic_vector( 5 downto 0);
    videoHSin_n : in std_logic;
    videoVSin_n : in std_logic;
    hCounterIn : in std_logic_vector(10 downto 0);
    vCounterIn : in std_logic_vector(10 downto 0);

    -- MODE
    PALMODE         : IN    STD_LOGIC;  -- caro
    interlaceMode : in std_logic;
    LEGACY_VGA      : IN    STD_LOGIC;
    
    -- Video Output
    videoRout : out std_logic_vector( 5 downto 0);
    videoGout : out std_logic_vector( 5 downto 0);
    videoBout : out std_logic_vector( 5 downto 0);
    videoHSout_n : out std_logic;
    videoVSout_n : out std_logic;
	BLANK_o         : OUT   STD_LOGIC;

	-- SWITCHED I/O SIGNALS
    RATIOMODE       : IN    STD_LOGIC_VECTOR( 2 DOWNTO 0)
    );
end vdp_vga;

architecture rtl of vdp_vga is
  -- video output enable
  signal videoOutX : std_logic;
--  signal videoOutY : std_logic;

  -- double buffer signal
  signal xPositionW : std_logic_vector(9 downto 0);
  signal xPositionR : std_logic_vector(9 downto 0);
  signal evenOdd    : std_logic;
  signal we_buf     : std_logic;
  signal dataRout   : std_logic_vector(5 downto 0);
  signal dataGout   : std_logic_vector(5 downto 0);
  signal dataBout   : std_logic_vector(5 downto 0);

  -- DISP_START_X + DISP_WIDTH < CLOCKS_PER_LINE/2 = 684
  constant DISP_WIDTH : integer := 562;  -- 30 + 512 + 20
  constant DISP_START_X : integer := 120;
begin

  videoRout <= dataRout when videoOutX = '1' else (others => '0');
  videoGout <= dataGout when videoOutX = '1' else (others => '0');
  videoBout <= dataBout when videoOutX = '1' else (others => '0');

  dbuf : work.VDP_DOUBLEBUF port map(clk21m, xPositionW, xPositionR, evenOdd, we_buf,
                            videoRin, videoGin, videoBin,
                            dataRout, dataGout, dataBout);

  xPositionW <= hCounterIn(10 downto 1) - (CLOCKS_PER_LINE/2 - DISP_WIDTH - 10);
  evenOdd <= vCounterIn(1);
  we_buf <= '1';
  
	BLANK_o <= '1' when VIDEOOUTX = '0' or FF_VSYNC_N = '0' else '0';

  process( clk21m, reset )
  begin
    if (reset = '1') then
      videoHSout_n <= '1';
      videoVSout_n <= '1';
      videoOutX <= '0';
      xPositionR <= (others => '0');
    elsif (clk21m'event and clk21m = '1') then

      -- Generate V-SYNC signal.
      -- The videoVSin_n signal is not used.
      if( interlaceMode = '0' ) then
        if( (vCounterIn = 3*2) or (vCounterIn = 524+3*2) )then
          videoVSout_n <= '0';
        elsif( (vCounterIn = 6*2) or (vCounterIn = 524+6*2) ) then
          videoVSout_n <= '1';
        end if;
      else
        if( (vCounterIn = 3*2) or (vCounterIn = 525+3*2) )then
          videoVSout_n <= '0';
        elsif( (vCounterIn = 6*2) or (vCounterIn = 525+6*2) ) then
          videoVSout_n <= '1';
        end if;
      end if;

      -- Generate H-SYNC signal.
      -- The videoHSin_n signal is not used.
      if( (hCounterIn = 0) or (hCounterIn = (CLOCKS_PER_LINE/2)) ) then
        videoHSout_n <= '0';
      elsif( (hCounterIn = 40) or (hCounterIn = (CLOCKS_PER_LINE/2) + 40) ) then
        videoHSout_n <= '1';
      end if;

      -- Generate data read timing.
      if( (hCounterIn = DISP_START_X) or
          (hCounterIn = DISP_START_X + (CLOCKS_PER_LINE/2)) ) then
        xPositionR <= (others => '0');
      else
        xPositionR <= xPositionR + 1;
      end if;

      -- Generate video output timing.
      if( (hCounterIn = DISP_START_X) or -- 120
          ((hCounterIn = DISP_START_X + (CLOCKS_PER_LINE/2)) and interlaceMode = '0') ) then
        videoOutX <= '1'; -- 120 a 682 or 804 to 1366 (if interlaced) 562 pixels total
      elsif( (hCounterIn = DISP_START_X+DISP_WIDTH) or -- 120 + 562 = 682
             (hCounterIn = DISP_START_X+DISP_WIDTH + (CLOCKS_PER_LINE/2)) ) then -- 120 + 562 + (1368/2) = 1366
				 
        videoOutX <= '0'; --out of the video area
      end if;
      
    end if;

  end process;
end rtl;




